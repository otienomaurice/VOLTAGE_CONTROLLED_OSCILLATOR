LTSpice Test Bench for V21
VCTRL vctrl 0 1
VRTN rtn 0 0
VFB vfb 0 5
VCAP vcap 0 2.5
VPOWER vpower 0 10
X1 rtn vcap vcc vctrl vfb  vlo vpower VCO_MauriceO
.options ITL1=1000
.DC VCTRL 0 5 0.1 VFB 0 5 5;* dc sweep
*.DC   VCTRL 0 5 0.1   VFB 0 5  5  VCAP 0.5 4.5 0.5
.include V21.sub
.end
